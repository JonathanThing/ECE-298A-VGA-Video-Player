/*
 * QSPI Module
 * Continuously reads 20-bit instructions from SPI flash
 */

 /* To Do: Rewrite with proper FSM format */

module qspi_controller (
    input  wire        clk,        // 25MHz pixel clock
    input  wire        rst_n,      // Reset (active low)
    
    // SPI Flash interface
    output wire        spi_clk,    // SPI clock = !clk
    output wire        spi_cs_n,   // Chip select (active low)
    output wire        spi_di,     // DI (data input to flash) - IO0
    output wire        spi_hold_n,   // HOLD (We have to hold it high during setup)

    input  wire        spi_io0,    // IO0 (for quad read)
    input  wire        spi_io1,     // DO (data output from flash) - IO1
    input  wire        spi_io2,    // IO2
    input  wire        spi_io3,     // IO3/HOLD

    input  wire        shift_data,  // Shift data through the buffers

    // Output interface
    output wire [17:0] instruction,        // 18-bit data output
    output wire        spi_cs_oe,
    output wire        spi_di_oe,
    output wire        spi_sclk_oe,
    output wire        spi_hold_n_oe,
    output wire        valid           // High when instruction is valid
);

    // State machine states
    localparam IDLE         = 3'b000;
    localparam SEND_CMD     = 3'b001;
    localparam DUMMY_CYCLES = 3'b010;
    localparam READ_DATA    = 3'b011;
    localparam WAIT_DATA    = 3'b111;

    // Internal signals
    reg [2:0]  state;
    reg [7:0]  bit_counter;
    reg [23:0] instruction_reg;
    reg        valid_reg;
    reg        cs_n_reg;
    reg        di_reg;
    reg [3:0]  oe_sig;      // 1 for output; 0 for input
    reg        hold_n_reg;
    reg        hold_read;
    
    wire [3:0] io_in_data;

    // SPI clock is inverted system clock
    assign spi_clk = !clk & !hold_read;
    assign spi_cs_n = cs_n_reg;
    assign spi_di = di_reg;
    assign spi_hold_n = hold_n_reg;

    // Quad data input (IO3, IO2, IO1/DO, IO0)
    assign io_in_data = {spi_io3, spi_io2, spi_io1, spi_io0};
    
    // Output assignments
    assign instruction = instruction_reg[17:0];
    assign valid = valid_reg;
    assign spi_cs_oe = oe_sig[0];
    assign spi_di_oe = oe_sig[1];
    assign spi_sclk_oe = oe_sig[2];
    assign spi_hold_n_oe = oe_sig[3];
    
    // Main state machine
    always @(posedge clk) begin
        if (!rst_n) begin
            state <= IDLE;
            bit_counter <= 8'b0;
            instruction_reg <= 24'b0;
            valid_reg <= 1'b0;
            cs_n_reg <= 1'b1;
            di_reg <= 1'b0;
            oe_sig <= 4'b0000;
            hold_n_reg <= 0;
        end else begin
            case (state)
                IDLE: begin
                    oe_sig <= 4'b1111;          
                    cs_n_reg <= 1'b1;          // Release chip select
                    bit_counter <= 8'b0;
                    valid_reg <= 1'b0;
                    di_reg <= 1'b0;
                    hold_n_reg <= 1;
                    hold_read <= 0;
                    state <= SEND_CMD;   
                end
                
                SEND_CMD: begin
                    cs_n_reg <= 1'b0;       // Pull CS low

                    // Send 8-bit command (6Bh = 01101011) on DI, MSB first
                    case (bit_counter)
                        0: di_reg <= 1'b0;  // bit 7
                        1: di_reg <= 1'b1;  // bit 6
                        2: di_reg <= 1'b1;  // bit 5
                        3: di_reg <= 1'b0;  // bit 4
                        4: di_reg <= 1'b1;  // bit 3
                        5: di_reg <= 1'b0;  // bit 2
                        6: di_reg <= 1'b1;  // bit 1
                        7: di_reg <= 1'b1;  // bit 0
                        default: di_reg <= 1'b0;
                    endcase
                    
                    bit_counter <= bit_counter + 1;

                    // We check 8 and not 7 because the SEND_CMD state starts one bit early
                    if (bit_counter == 8) begin  
                        state <= DUMMY_CYCLES;
                        bit_counter <= 8'b0;
                    end
                end
                
                DUMMY_CYCLES: begin
                    // Wait for dummy cycles (32 dummy clocks as per datasheet)
                    di_reg <= 1'b0;  // Keep DI low during dummy cycles
                    bit_counter <= bit_counter + 1;

                    if (bit_counter == 31) begin  // 31 cycles already occured,
                        oe_sig <= 4'b0101;
                        state <= READ_DATA;
                        bit_counter <= 8'b0;
                    end
                end
                
                READ_DATA: begin
                    
                    // Read 24 bits of data (6 cycles of 4 bits each)
                    instruction_reg <= {instruction_reg[19:0], io_in_data};
                    bit_counter <= bit_counter + 1;
                    
                    if (bit_counter == 5) begin  // 3 bytes received (6 cycles)
                        valid_reg <= 1'b1;
                        bit_counter <= 8'b0;
                        if (!shift_data) begin
                            state <= WAIT_DATA;
                        end
                    end else begin
                        valid_reg <= 1'b0;
                    end
                end

                WAIT_DATA: begin        
                    hold_read <= 1'b1;
                    if (shift_data) begin   // Wait for data to be consumed until reading next message
                        state <= READ_DATA;
                        hold_read <= 1'b0;
                        bit_counter <= 8'b0;
                    end
                end

                default: begin
                    state <= IDLE;
                    oe_sig <= 4'b1101;
                    hold_n_reg <= 0;
                end
            endcase
        end
    end

endmodule